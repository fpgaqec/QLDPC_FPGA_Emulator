library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.LLR_fpQLP127x254_q_pkg.all;

package LLR_fpQLP127x254_q_em_pkg is
	--generics
	constant Ng: integer:= 40; -- #png 
	constant Mg: integer:= 7; -- #clock cycles S/P 
	constant Nvnu: integer:= 254; -- #VNUs  
	constant M_Hlogic: integer:= 14; -- #M_Hlogic  
	constant M_buf: integer:= 8; -- #Buffer words   
	constant A_buf: integer:= 3; -- #Buffer address bus  
	constant N_ram: integer:= 512; -- #words RAM  
	constant A_ram: integer:= 9;  -- #bits RAM address  
	constant ESC_DLOOP_CNT: integer:= 0;  -- Scaling read Dloop_cnt  
	--generic for implementation/simpulation
	constant DEBUG: integer := 1; -- Debug mode 
	--generics for simpulation
	constant Mloop: integer:= 31; -- #iterations  
	constant Nerrors: integer:= 1; -- #errors  
	constant Threshold: integer:= -14342; -- #threshold  

	--TB signals
	signal db_cmp_s : std_logic_vector(0 to Ng-1); 
	signal db_run : std_logic; 
	signal db_load : std_logic; 
	signal db_b1_edec_s : std_logic; 
	signal db_b7_edec_r : std_logic; 
	signal db_b8_edec_r : std_logic; 
	signal db_b9_edec_r : std_logic; 
	signal db_llr_block : p_type_a254xQIstd; 
	signal db_b4_dec_block_s: std_logic_vector(0 to 253); 
	signal db_b4_parity_check_r : std_logic; 
	signal db_b8_errf_cnt_r : unsigned(15 downto 0); 
	signal db_b8_errl_cnt_r : unsigned(15 downto 0); 
	signal db_b9_dloop_cnt_r : unsigned(85 downto 0); 
	signal db_b7_dec_cnt_r: unsigned(79 downto 0); 

	--types

	--constraints
	constant cnt_llr_in: p_type_a254xQIstd := ("1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000",
	                                           "1111000");

--
end package;
