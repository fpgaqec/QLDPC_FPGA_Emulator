library ieee;
use ieee.std_logic_1164.all;
use work.LLR_fpQLP127x254_q_pkg.all;

entity LLR_fpQLP127x254_xH is 
	port(id_noixe_block : in std_logic_vector(0 to 253); -- noisex : 1 bit 
	     od_syn_block : out p_type_a127xstd); -- syndrome block : 1 bit
end LLR_fpQLP127x254_xH; 
 
architecture rtl of LLR_fpQLP127x254_xH is 
begin 
	od_syn_block(0) <= id_noixe_block(0) xor id_noixe_block(18) xor id_noixe_block(53) xor id_noixe_block(127) xor id_noixe_block(139) xor id_noixe_block(252);
	od_syn_block(1) <= id_noixe_block(1) xor id_noixe_block(19) xor id_noixe_block(54) xor id_noixe_block(128) xor id_noixe_block(140) xor id_noixe_block(253);
	od_syn_block(2) <= id_noixe_block(2) xor id_noixe_block(20) xor id_noixe_block(55) xor id_noixe_block(127) xor id_noixe_block(129) xor id_noixe_block(141);
	od_syn_block(3) <= id_noixe_block(3) xor id_noixe_block(21) xor id_noixe_block(56) xor id_noixe_block(128) xor id_noixe_block(130) xor id_noixe_block(142);
	od_syn_block(4) <= id_noixe_block(4) xor id_noixe_block(22) xor id_noixe_block(57) xor id_noixe_block(129) xor id_noixe_block(131) xor id_noixe_block(143);
	od_syn_block(5) <= id_noixe_block(5) xor id_noixe_block(23) xor id_noixe_block(58) xor id_noixe_block(130) xor id_noixe_block(132) xor id_noixe_block(144);
	od_syn_block(6) <= id_noixe_block(6) xor id_noixe_block(24) xor id_noixe_block(59) xor id_noixe_block(131) xor id_noixe_block(133) xor id_noixe_block(145);
	od_syn_block(7) <= id_noixe_block(7) xor id_noixe_block(25) xor id_noixe_block(60) xor id_noixe_block(132) xor id_noixe_block(134) xor id_noixe_block(146);
	od_syn_block(8) <= id_noixe_block(8) xor id_noixe_block(26) xor id_noixe_block(61) xor id_noixe_block(133) xor id_noixe_block(135) xor id_noixe_block(147);
	od_syn_block(9) <= id_noixe_block(9) xor id_noixe_block(27) xor id_noixe_block(62) xor id_noixe_block(134) xor id_noixe_block(136) xor id_noixe_block(148);
	od_syn_block(10) <= id_noixe_block(10) xor id_noixe_block(28) xor id_noixe_block(63) xor id_noixe_block(135) xor id_noixe_block(137) xor id_noixe_block(149);
	od_syn_block(11) <= id_noixe_block(11) xor id_noixe_block(29) xor id_noixe_block(64) xor id_noixe_block(136) xor id_noixe_block(138) xor id_noixe_block(150);
	od_syn_block(12) <= id_noixe_block(12) xor id_noixe_block(30) xor id_noixe_block(65) xor id_noixe_block(137) xor id_noixe_block(139) xor id_noixe_block(151);
	od_syn_block(13) <= id_noixe_block(13) xor id_noixe_block(31) xor id_noixe_block(66) xor id_noixe_block(138) xor id_noixe_block(140) xor id_noixe_block(152);
	od_syn_block(14) <= id_noixe_block(14) xor id_noixe_block(32) xor id_noixe_block(67) xor id_noixe_block(139) xor id_noixe_block(141) xor id_noixe_block(153);
	od_syn_block(15) <= id_noixe_block(15) xor id_noixe_block(33) xor id_noixe_block(68) xor id_noixe_block(140) xor id_noixe_block(142) xor id_noixe_block(154);
	od_syn_block(16) <= id_noixe_block(16) xor id_noixe_block(34) xor id_noixe_block(69) xor id_noixe_block(141) xor id_noixe_block(143) xor id_noixe_block(155);
	od_syn_block(17) <= id_noixe_block(17) xor id_noixe_block(35) xor id_noixe_block(70) xor id_noixe_block(142) xor id_noixe_block(144) xor id_noixe_block(156);
	od_syn_block(18) <= id_noixe_block(18) xor id_noixe_block(36) xor id_noixe_block(71) xor id_noixe_block(143) xor id_noixe_block(145) xor id_noixe_block(157);
	od_syn_block(19) <= id_noixe_block(19) xor id_noixe_block(37) xor id_noixe_block(72) xor id_noixe_block(144) xor id_noixe_block(146) xor id_noixe_block(158);
	od_syn_block(20) <= id_noixe_block(20) xor id_noixe_block(38) xor id_noixe_block(73) xor id_noixe_block(145) xor id_noixe_block(147) xor id_noixe_block(159);
	od_syn_block(21) <= id_noixe_block(21) xor id_noixe_block(39) xor id_noixe_block(74) xor id_noixe_block(146) xor id_noixe_block(148) xor id_noixe_block(160);
	od_syn_block(22) <= id_noixe_block(22) xor id_noixe_block(40) xor id_noixe_block(75) xor id_noixe_block(147) xor id_noixe_block(149) xor id_noixe_block(161);
	od_syn_block(23) <= id_noixe_block(23) xor id_noixe_block(41) xor id_noixe_block(76) xor id_noixe_block(148) xor id_noixe_block(150) xor id_noixe_block(162);
	od_syn_block(24) <= id_noixe_block(24) xor id_noixe_block(42) xor id_noixe_block(77) xor id_noixe_block(149) xor id_noixe_block(151) xor id_noixe_block(163);
	od_syn_block(25) <= id_noixe_block(25) xor id_noixe_block(43) xor id_noixe_block(78) xor id_noixe_block(150) xor id_noixe_block(152) xor id_noixe_block(164);
	od_syn_block(26) <= id_noixe_block(26) xor id_noixe_block(44) xor id_noixe_block(79) xor id_noixe_block(151) xor id_noixe_block(153) xor id_noixe_block(165);
	od_syn_block(27) <= id_noixe_block(27) xor id_noixe_block(45) xor id_noixe_block(80) xor id_noixe_block(152) xor id_noixe_block(154) xor id_noixe_block(166);
	od_syn_block(28) <= id_noixe_block(28) xor id_noixe_block(46) xor id_noixe_block(81) xor id_noixe_block(153) xor id_noixe_block(155) xor id_noixe_block(167);
	od_syn_block(29) <= id_noixe_block(29) xor id_noixe_block(47) xor id_noixe_block(82) xor id_noixe_block(154) xor id_noixe_block(156) xor id_noixe_block(168);
	od_syn_block(30) <= id_noixe_block(30) xor id_noixe_block(48) xor id_noixe_block(83) xor id_noixe_block(155) xor id_noixe_block(157) xor id_noixe_block(169);
	od_syn_block(31) <= id_noixe_block(31) xor id_noixe_block(49) xor id_noixe_block(84) xor id_noixe_block(156) xor id_noixe_block(158) xor id_noixe_block(170);
	od_syn_block(32) <= id_noixe_block(32) xor id_noixe_block(50) xor id_noixe_block(85) xor id_noixe_block(157) xor id_noixe_block(159) xor id_noixe_block(171);
	od_syn_block(33) <= id_noixe_block(33) xor id_noixe_block(51) xor id_noixe_block(86) xor id_noixe_block(158) xor id_noixe_block(160) xor id_noixe_block(172);
	od_syn_block(34) <= id_noixe_block(34) xor id_noixe_block(52) xor id_noixe_block(87) xor id_noixe_block(159) xor id_noixe_block(161) xor id_noixe_block(173);
	od_syn_block(35) <= id_noixe_block(35) xor id_noixe_block(53) xor id_noixe_block(88) xor id_noixe_block(160) xor id_noixe_block(162) xor id_noixe_block(174);
	od_syn_block(36) <= id_noixe_block(36) xor id_noixe_block(54) xor id_noixe_block(89) xor id_noixe_block(161) xor id_noixe_block(163) xor id_noixe_block(175);
	od_syn_block(37) <= id_noixe_block(37) xor id_noixe_block(55) xor id_noixe_block(90) xor id_noixe_block(162) xor id_noixe_block(164) xor id_noixe_block(176);
	od_syn_block(38) <= id_noixe_block(38) xor id_noixe_block(56) xor id_noixe_block(91) xor id_noixe_block(163) xor id_noixe_block(165) xor id_noixe_block(177);
	od_syn_block(39) <= id_noixe_block(39) xor id_noixe_block(57) xor id_noixe_block(92) xor id_noixe_block(164) xor id_noixe_block(166) xor id_noixe_block(178);
	od_syn_block(40) <= id_noixe_block(40) xor id_noixe_block(58) xor id_noixe_block(93) xor id_noixe_block(165) xor id_noixe_block(167) xor id_noixe_block(179);
	od_syn_block(41) <= id_noixe_block(41) xor id_noixe_block(59) xor id_noixe_block(94) xor id_noixe_block(166) xor id_noixe_block(168) xor id_noixe_block(180);
	od_syn_block(42) <= id_noixe_block(42) xor id_noixe_block(60) xor id_noixe_block(95) xor id_noixe_block(167) xor id_noixe_block(169) xor id_noixe_block(181);
	od_syn_block(43) <= id_noixe_block(43) xor id_noixe_block(61) xor id_noixe_block(96) xor id_noixe_block(168) xor id_noixe_block(170) xor id_noixe_block(182);
	od_syn_block(44) <= id_noixe_block(44) xor id_noixe_block(62) xor id_noixe_block(97) xor id_noixe_block(169) xor id_noixe_block(171) xor id_noixe_block(183);
	od_syn_block(45) <= id_noixe_block(45) xor id_noixe_block(63) xor id_noixe_block(98) xor id_noixe_block(170) xor id_noixe_block(172) xor id_noixe_block(184);
	od_syn_block(46) <= id_noixe_block(46) xor id_noixe_block(64) xor id_noixe_block(99) xor id_noixe_block(171) xor id_noixe_block(173) xor id_noixe_block(185);
	od_syn_block(47) <= id_noixe_block(47) xor id_noixe_block(65) xor id_noixe_block(100) xor id_noixe_block(172) xor id_noixe_block(174) xor id_noixe_block(186);
	od_syn_block(48) <= id_noixe_block(48) xor id_noixe_block(66) xor id_noixe_block(101) xor id_noixe_block(173) xor id_noixe_block(175) xor id_noixe_block(187);
	od_syn_block(49) <= id_noixe_block(49) xor id_noixe_block(67) xor id_noixe_block(102) xor id_noixe_block(174) xor id_noixe_block(176) xor id_noixe_block(188);
	od_syn_block(50) <= id_noixe_block(50) xor id_noixe_block(68) xor id_noixe_block(103) xor id_noixe_block(175) xor id_noixe_block(177) xor id_noixe_block(189);
	od_syn_block(51) <= id_noixe_block(51) xor id_noixe_block(69) xor id_noixe_block(104) xor id_noixe_block(176) xor id_noixe_block(178) xor id_noixe_block(190);
	od_syn_block(52) <= id_noixe_block(52) xor id_noixe_block(70) xor id_noixe_block(105) xor id_noixe_block(177) xor id_noixe_block(179) xor id_noixe_block(191);
	od_syn_block(53) <= id_noixe_block(53) xor id_noixe_block(71) xor id_noixe_block(106) xor id_noixe_block(178) xor id_noixe_block(180) xor id_noixe_block(192);
	od_syn_block(54) <= id_noixe_block(54) xor id_noixe_block(72) xor id_noixe_block(107) xor id_noixe_block(179) xor id_noixe_block(181) xor id_noixe_block(193);
	od_syn_block(55) <= id_noixe_block(55) xor id_noixe_block(73) xor id_noixe_block(108) xor id_noixe_block(180) xor id_noixe_block(182) xor id_noixe_block(194);
	od_syn_block(56) <= id_noixe_block(56) xor id_noixe_block(74) xor id_noixe_block(109) xor id_noixe_block(181) xor id_noixe_block(183) xor id_noixe_block(195);
	od_syn_block(57) <= id_noixe_block(57) xor id_noixe_block(75) xor id_noixe_block(110) xor id_noixe_block(182) xor id_noixe_block(184) xor id_noixe_block(196);
	od_syn_block(58) <= id_noixe_block(58) xor id_noixe_block(76) xor id_noixe_block(111) xor id_noixe_block(183) xor id_noixe_block(185) xor id_noixe_block(197);
	od_syn_block(59) <= id_noixe_block(59) xor id_noixe_block(77) xor id_noixe_block(112) xor id_noixe_block(184) xor id_noixe_block(186) xor id_noixe_block(198);
	od_syn_block(60) <= id_noixe_block(60) xor id_noixe_block(78) xor id_noixe_block(113) xor id_noixe_block(185) xor id_noixe_block(187) xor id_noixe_block(199);
	od_syn_block(61) <= id_noixe_block(61) xor id_noixe_block(79) xor id_noixe_block(114) xor id_noixe_block(186) xor id_noixe_block(188) xor id_noixe_block(200);
	od_syn_block(62) <= id_noixe_block(62) xor id_noixe_block(80) xor id_noixe_block(115) xor id_noixe_block(187) xor id_noixe_block(189) xor id_noixe_block(201);
	od_syn_block(63) <= id_noixe_block(63) xor id_noixe_block(81) xor id_noixe_block(116) xor id_noixe_block(188) xor id_noixe_block(190) xor id_noixe_block(202);
	od_syn_block(64) <= id_noixe_block(64) xor id_noixe_block(82) xor id_noixe_block(117) xor id_noixe_block(189) xor id_noixe_block(191) xor id_noixe_block(203);
	od_syn_block(65) <= id_noixe_block(65) xor id_noixe_block(83) xor id_noixe_block(118) xor id_noixe_block(190) xor id_noixe_block(192) xor id_noixe_block(204);
	od_syn_block(66) <= id_noixe_block(66) xor id_noixe_block(84) xor id_noixe_block(119) xor id_noixe_block(191) xor id_noixe_block(193) xor id_noixe_block(205);
	od_syn_block(67) <= id_noixe_block(67) xor id_noixe_block(85) xor id_noixe_block(120) xor id_noixe_block(192) xor id_noixe_block(194) xor id_noixe_block(206);
	od_syn_block(68) <= id_noixe_block(68) xor id_noixe_block(86) xor id_noixe_block(121) xor id_noixe_block(193) xor id_noixe_block(195) xor id_noixe_block(207);
	od_syn_block(69) <= id_noixe_block(69) xor id_noixe_block(87) xor id_noixe_block(122) xor id_noixe_block(194) xor id_noixe_block(196) xor id_noixe_block(208);
	od_syn_block(70) <= id_noixe_block(70) xor id_noixe_block(88) xor id_noixe_block(123) xor id_noixe_block(195) xor id_noixe_block(197) xor id_noixe_block(209);
	od_syn_block(71) <= id_noixe_block(71) xor id_noixe_block(89) xor id_noixe_block(124) xor id_noixe_block(196) xor id_noixe_block(198) xor id_noixe_block(210);
	od_syn_block(72) <= id_noixe_block(72) xor id_noixe_block(90) xor id_noixe_block(125) xor id_noixe_block(197) xor id_noixe_block(199) xor id_noixe_block(211);
	od_syn_block(73) <= id_noixe_block(73) xor id_noixe_block(91) xor id_noixe_block(126) xor id_noixe_block(198) xor id_noixe_block(200) xor id_noixe_block(212);
	od_syn_block(74) <= id_noixe_block(0) xor id_noixe_block(74) xor id_noixe_block(92) xor id_noixe_block(199) xor id_noixe_block(201) xor id_noixe_block(213);
	od_syn_block(75) <= id_noixe_block(1) xor id_noixe_block(75) xor id_noixe_block(93) xor id_noixe_block(200) xor id_noixe_block(202) xor id_noixe_block(214);
	od_syn_block(76) <= id_noixe_block(2) xor id_noixe_block(76) xor id_noixe_block(94) xor id_noixe_block(201) xor id_noixe_block(203) xor id_noixe_block(215);
	od_syn_block(77) <= id_noixe_block(3) xor id_noixe_block(77) xor id_noixe_block(95) xor id_noixe_block(202) xor id_noixe_block(204) xor id_noixe_block(216);
	od_syn_block(78) <= id_noixe_block(4) xor id_noixe_block(78) xor id_noixe_block(96) xor id_noixe_block(203) xor id_noixe_block(205) xor id_noixe_block(217);
	od_syn_block(79) <= id_noixe_block(5) xor id_noixe_block(79) xor id_noixe_block(97) xor id_noixe_block(204) xor id_noixe_block(206) xor id_noixe_block(218);
	od_syn_block(80) <= id_noixe_block(6) xor id_noixe_block(80) xor id_noixe_block(98) xor id_noixe_block(205) xor id_noixe_block(207) xor id_noixe_block(219);
	od_syn_block(81) <= id_noixe_block(7) xor id_noixe_block(81) xor id_noixe_block(99) xor id_noixe_block(206) xor id_noixe_block(208) xor id_noixe_block(220);
	od_syn_block(82) <= id_noixe_block(8) xor id_noixe_block(82) xor id_noixe_block(100) xor id_noixe_block(207) xor id_noixe_block(209) xor id_noixe_block(221);
	od_syn_block(83) <= id_noixe_block(9) xor id_noixe_block(83) xor id_noixe_block(101) xor id_noixe_block(208) xor id_noixe_block(210) xor id_noixe_block(222);
	od_syn_block(84) <= id_noixe_block(10) xor id_noixe_block(84) xor id_noixe_block(102) xor id_noixe_block(209) xor id_noixe_block(211) xor id_noixe_block(223);
	od_syn_block(85) <= id_noixe_block(11) xor id_noixe_block(85) xor id_noixe_block(103) xor id_noixe_block(210) xor id_noixe_block(212) xor id_noixe_block(224);
	od_syn_block(86) <= id_noixe_block(12) xor id_noixe_block(86) xor id_noixe_block(104) xor id_noixe_block(211) xor id_noixe_block(213) xor id_noixe_block(225);
	od_syn_block(87) <= id_noixe_block(13) xor id_noixe_block(87) xor id_noixe_block(105) xor id_noixe_block(212) xor id_noixe_block(214) xor id_noixe_block(226);
	od_syn_block(88) <= id_noixe_block(14) xor id_noixe_block(88) xor id_noixe_block(106) xor id_noixe_block(213) xor id_noixe_block(215) xor id_noixe_block(227);
	od_syn_block(89) <= id_noixe_block(15) xor id_noixe_block(89) xor id_noixe_block(107) xor id_noixe_block(214) xor id_noixe_block(216) xor id_noixe_block(228);
	od_syn_block(90) <= id_noixe_block(16) xor id_noixe_block(90) xor id_noixe_block(108) xor id_noixe_block(215) xor id_noixe_block(217) xor id_noixe_block(229);
	od_syn_block(91) <= id_noixe_block(17) xor id_noixe_block(91) xor id_noixe_block(109) xor id_noixe_block(216) xor id_noixe_block(218) xor id_noixe_block(230);
	od_syn_block(92) <= id_noixe_block(18) xor id_noixe_block(92) xor id_noixe_block(110) xor id_noixe_block(217) xor id_noixe_block(219) xor id_noixe_block(231);
	od_syn_block(93) <= id_noixe_block(19) xor id_noixe_block(93) xor id_noixe_block(111) xor id_noixe_block(218) xor id_noixe_block(220) xor id_noixe_block(232);
	od_syn_block(94) <= id_noixe_block(20) xor id_noixe_block(94) xor id_noixe_block(112) xor id_noixe_block(219) xor id_noixe_block(221) xor id_noixe_block(233);
	od_syn_block(95) <= id_noixe_block(21) xor id_noixe_block(95) xor id_noixe_block(113) xor id_noixe_block(220) xor id_noixe_block(222) xor id_noixe_block(234);
	od_syn_block(96) <= id_noixe_block(22) xor id_noixe_block(96) xor id_noixe_block(114) xor id_noixe_block(221) xor id_noixe_block(223) xor id_noixe_block(235);
	od_syn_block(97) <= id_noixe_block(23) xor id_noixe_block(97) xor id_noixe_block(115) xor id_noixe_block(222) xor id_noixe_block(224) xor id_noixe_block(236);
	od_syn_block(98) <= id_noixe_block(24) xor id_noixe_block(98) xor id_noixe_block(116) xor id_noixe_block(223) xor id_noixe_block(225) xor id_noixe_block(237);
	od_syn_block(99) <= id_noixe_block(25) xor id_noixe_block(99) xor id_noixe_block(117) xor id_noixe_block(224) xor id_noixe_block(226) xor id_noixe_block(238);
	od_syn_block(100) <= id_noixe_block(26) xor id_noixe_block(100) xor id_noixe_block(118) xor id_noixe_block(225) xor id_noixe_block(227) xor id_noixe_block(239);
	od_syn_block(101) <= id_noixe_block(27) xor id_noixe_block(101) xor id_noixe_block(119) xor id_noixe_block(226) xor id_noixe_block(228) xor id_noixe_block(240);
	od_syn_block(102) <= id_noixe_block(28) xor id_noixe_block(102) xor id_noixe_block(120) xor id_noixe_block(227) xor id_noixe_block(229) xor id_noixe_block(241);
	od_syn_block(103) <= id_noixe_block(29) xor id_noixe_block(103) xor id_noixe_block(121) xor id_noixe_block(228) xor id_noixe_block(230) xor id_noixe_block(242);
	od_syn_block(104) <= id_noixe_block(30) xor id_noixe_block(104) xor id_noixe_block(122) xor id_noixe_block(229) xor id_noixe_block(231) xor id_noixe_block(243);
	od_syn_block(105) <= id_noixe_block(31) xor id_noixe_block(105) xor id_noixe_block(123) xor id_noixe_block(230) xor id_noixe_block(232) xor id_noixe_block(244);
	od_syn_block(106) <= id_noixe_block(32) xor id_noixe_block(106) xor id_noixe_block(124) xor id_noixe_block(231) xor id_noixe_block(233) xor id_noixe_block(245);
	od_syn_block(107) <= id_noixe_block(33) xor id_noixe_block(107) xor id_noixe_block(125) xor id_noixe_block(232) xor id_noixe_block(234) xor id_noixe_block(246);
	od_syn_block(108) <= id_noixe_block(34) xor id_noixe_block(108) xor id_noixe_block(126) xor id_noixe_block(233) xor id_noixe_block(235) xor id_noixe_block(247);
	od_syn_block(109) <= id_noixe_block(0) xor id_noixe_block(35) xor id_noixe_block(109) xor id_noixe_block(234) xor id_noixe_block(236) xor id_noixe_block(248);
	od_syn_block(110) <= id_noixe_block(1) xor id_noixe_block(36) xor id_noixe_block(110) xor id_noixe_block(235) xor id_noixe_block(237) xor id_noixe_block(249);
	od_syn_block(111) <= id_noixe_block(2) xor id_noixe_block(37) xor id_noixe_block(111) xor id_noixe_block(236) xor id_noixe_block(238) xor id_noixe_block(250);
	od_syn_block(112) <= id_noixe_block(3) xor id_noixe_block(38) xor id_noixe_block(112) xor id_noixe_block(237) xor id_noixe_block(239) xor id_noixe_block(251);
	od_syn_block(113) <= id_noixe_block(4) xor id_noixe_block(39) xor id_noixe_block(113) xor id_noixe_block(238) xor id_noixe_block(240) xor id_noixe_block(252);
	od_syn_block(114) <= id_noixe_block(5) xor id_noixe_block(40) xor id_noixe_block(114) xor id_noixe_block(239) xor id_noixe_block(241) xor id_noixe_block(253);
	od_syn_block(115) <= id_noixe_block(6) xor id_noixe_block(41) xor id_noixe_block(115) xor id_noixe_block(127) xor id_noixe_block(240) xor id_noixe_block(242);
	od_syn_block(116) <= id_noixe_block(7) xor id_noixe_block(42) xor id_noixe_block(116) xor id_noixe_block(128) xor id_noixe_block(241) xor id_noixe_block(243);
	od_syn_block(117) <= id_noixe_block(8) xor id_noixe_block(43) xor id_noixe_block(117) xor id_noixe_block(129) xor id_noixe_block(242) xor id_noixe_block(244);
	od_syn_block(118) <= id_noixe_block(9) xor id_noixe_block(44) xor id_noixe_block(118) xor id_noixe_block(130) xor id_noixe_block(243) xor id_noixe_block(245);
	od_syn_block(119) <= id_noixe_block(10) xor id_noixe_block(45) xor id_noixe_block(119) xor id_noixe_block(131) xor id_noixe_block(244) xor id_noixe_block(246);
	od_syn_block(120) <= id_noixe_block(11) xor id_noixe_block(46) xor id_noixe_block(120) xor id_noixe_block(132) xor id_noixe_block(245) xor id_noixe_block(247);
	od_syn_block(121) <= id_noixe_block(12) xor id_noixe_block(47) xor id_noixe_block(121) xor id_noixe_block(133) xor id_noixe_block(246) xor id_noixe_block(248);
	od_syn_block(122) <= id_noixe_block(13) xor id_noixe_block(48) xor id_noixe_block(122) xor id_noixe_block(134) xor id_noixe_block(247) xor id_noixe_block(249);
	od_syn_block(123) <= id_noixe_block(14) xor id_noixe_block(49) xor id_noixe_block(123) xor id_noixe_block(135) xor id_noixe_block(248) xor id_noixe_block(250);
	od_syn_block(124) <= id_noixe_block(15) xor id_noixe_block(50) xor id_noixe_block(124) xor id_noixe_block(136) xor id_noixe_block(249) xor id_noixe_block(251);
	od_syn_block(125) <= id_noixe_block(16) xor id_noixe_block(51) xor id_noixe_block(125) xor id_noixe_block(137) xor id_noixe_block(250) xor id_noixe_block(252);
	od_syn_block(126) <= id_noixe_block(17) xor id_noixe_block(52) xor id_noixe_block(126) xor id_noixe_block(138) xor id_noixe_block(251) xor id_noixe_block(253);
end rtl; 
