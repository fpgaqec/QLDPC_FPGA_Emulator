library ieee;
use ieee.std_logic_1164.all;
use work.LLR_fpQLP127x254_q_pkg.all;

entity LLR_fpQLP127x254_xHlogic is 
	port(id_xor_block : in std_logic_vector(0 to 253); -- check xor : 1 bit 
	     od_logic_block : out std_logic_vector(0 to 13)); -- logic : 1 bit 
end LLR_fpQLP127x254_xHlogic; 
 
architecture rtl of LLR_fpQLP127x254_xHlogic is 
begin 
	od_logic_block(0) <= id_xor_block(120) xor id_xor_block(121) xor id_xor_block(122) xor id_xor_block(123) xor id_xor_block(124) xor id_xor_block(125) xor id_xor_block(126) xor id_xor_block(129) xor id_xor_block(130) xor id_xor_block(133) xor id_xor_block(134) xor id_xor_block(135) xor id_xor_block(136) xor id_xor_block(139) xor id_xor_block(140) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(143) xor id_xor_block(144) xor id_xor_block(145) xor id_xor_block(148) xor id_xor_block(149) xor id_xor_block(150) xor id_xor_block(154) xor id_xor_block(155) xor id_xor_block(156) xor id_xor_block(164) xor id_xor_block(165) xor id_xor_block(167) xor id_xor_block(168) xor id_xor_block(172) xor id_xor_block(173) xor id_xor_block(174) xor id_xor_block(185) xor id_xor_block(187) xor id_xor_block(188) xor id_xor_block(189) xor id_xor_block(190) xor id_xor_block(191) xor id_xor_block(193) xor id_xor_block(194) xor id_xor_block(195) xor id_xor_block(196) xor id_xor_block(197) xor id_xor_block(198) xor id_xor_block(201) xor id_xor_block(202) xor id_xor_block(205) xor id_xor_block(206) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(214) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(217) xor id_xor_block(218) xor id_xor_block(219) xor id_xor_block(221) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(225) xor id_xor_block(226) xor id_xor_block(227) xor id_xor_block(229) xor id_xor_block(230) xor id_xor_block(231) xor id_xor_block(232) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(235) xor id_xor_block(236) xor id_xor_block(237) xor id_xor_block(238) xor id_xor_block(239) xor id_xor_block(240);
	od_logic_block(1) <= id_xor_block(120) xor id_xor_block(126) xor id_xor_block(127) xor id_xor_block(129) xor id_xor_block(131) xor id_xor_block(133) xor id_xor_block(137) xor id_xor_block(139) xor id_xor_block(142) xor id_xor_block(143) xor id_xor_block(145) xor id_xor_block(146) xor id_xor_block(148) xor id_xor_block(151) xor id_xor_block(154) xor id_xor_block(157) xor id_xor_block(159) xor id_xor_block(160) xor id_xor_block(163) xor id_xor_block(164) xor id_xor_block(166) xor id_xor_block(167) xor id_xor_block(169) xor id_xor_block(172) xor id_xor_block(175) xor id_xor_block(177) xor id_xor_block(178) xor id_xor_block(180) xor id_xor_block(181) xor id_xor_block(185) xor id_xor_block(186) xor id_xor_block(187) xor id_xor_block(192) xor id_xor_block(193) xor id_xor_block(201) xor id_xor_block(203) xor id_xor_block(205) xor id_xor_block(207) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(216) xor id_xor_block(217) xor id_xor_block(220) xor id_xor_block(221) xor id_xor_block(222) xor id_xor_block(223) xor id_xor_block(228) xor id_xor_block(229) xor id_xor_block(233) xor id_xor_block(235) xor id_xor_block(241);
	od_logic_block(2) <= id_xor_block(121) xor id_xor_block(126) xor id_xor_block(127) xor id_xor_block(128) xor id_xor_block(130) xor id_xor_block(132) xor id_xor_block(134) xor id_xor_block(138) xor id_xor_block(140) xor id_xor_block(142) xor id_xor_block(144) xor id_xor_block(145) xor id_xor_block(146) xor id_xor_block(147) xor id_xor_block(149) xor id_xor_block(152) xor id_xor_block(155) xor id_xor_block(158) xor id_xor_block(159) xor id_xor_block(161) xor id_xor_block(163) xor id_xor_block(164) xor id_xor_block(165) xor id_xor_block(167) xor id_xor_block(168) xor id_xor_block(170) xor id_xor_block(173) xor id_xor_block(176) xor id_xor_block(177) xor id_xor_block(179) xor id_xor_block(180) xor id_xor_block(182) xor id_xor_block(186) xor id_xor_block(187) xor id_xor_block(188) xor id_xor_block(193) xor id_xor_block(194) xor id_xor_block(199) xor id_xor_block(202) xor id_xor_block(204) xor id_xor_block(206) xor id_xor_block(208) xor id_xor_block(214) xor id_xor_block(216) xor id_xor_block(218) xor id_xor_block(221) xor id_xor_block(222) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(229) xor id_xor_block(230) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(235) xor id_xor_block(236) xor id_xor_block(242);
	od_logic_block(3) <= id_xor_block(122) xor id_xor_block(126) xor id_xor_block(127) xor id_xor_block(128) xor id_xor_block(129) xor id_xor_block(131) xor id_xor_block(133) xor id_xor_block(135) xor id_xor_block(139) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(146) xor id_xor_block(147) xor id_xor_block(148) xor id_xor_block(150) xor id_xor_block(153) xor id_xor_block(156) xor id_xor_block(162) xor id_xor_block(163) xor id_xor_block(164) xor id_xor_block(165) xor id_xor_block(166) xor id_xor_block(168) xor id_xor_block(169) xor id_xor_block(171) xor id_xor_block(174) xor id_xor_block(183) xor id_xor_block(187) xor id_xor_block(188) xor id_xor_block(189) xor id_xor_block(194) xor id_xor_block(195) xor id_xor_block(199) xor id_xor_block(200) xor id_xor_block(203) xor id_xor_block(205) xor id_xor_block(207) xor id_xor_block(209) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(219) xor id_xor_block(222) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(225) xor id_xor_block(230) xor id_xor_block(231) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(236) xor id_xor_block(237) xor id_xor_block(243);
	od_logic_block(4) <= id_xor_block(123) xor id_xor_block(126) xor id_xor_block(127) xor id_xor_block(128) xor id_xor_block(129) xor id_xor_block(130) xor id_xor_block(132) xor id_xor_block(134) xor id_xor_block(136) xor id_xor_block(140) xor id_xor_block(145) xor id_xor_block(147) xor id_xor_block(148) xor id_xor_block(149) xor id_xor_block(151) xor id_xor_block(154) xor id_xor_block(157) xor id_xor_block(159) xor id_xor_block(160) xor id_xor_block(164) xor id_xor_block(165) xor id_xor_block(166) xor id_xor_block(167) xor id_xor_block(169) xor id_xor_block(170) xor id_xor_block(172) xor id_xor_block(175) xor id_xor_block(177) xor id_xor_block(178) xor id_xor_block(180) xor id_xor_block(181) xor id_xor_block(184) xor id_xor_block(188) xor id_xor_block(189) xor id_xor_block(190) xor id_xor_block(195) xor id_xor_block(196) xor id_xor_block(199) xor id_xor_block(200) xor id_xor_block(201) xor id_xor_block(204) xor id_xor_block(206) xor id_xor_block(208) xor id_xor_block(210) xor id_xor_block(212) xor id_xor_block(214) xor id_xor_block(220) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(225) xor id_xor_block(226) xor id_xor_block(231) xor id_xor_block(232) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(237) xor id_xor_block(238) xor id_xor_block(244);
	od_logic_block(5) <= id_xor_block(124) xor id_xor_block(126) xor id_xor_block(127) xor id_xor_block(128) xor id_xor_block(129) xor id_xor_block(130) xor id_xor_block(131) xor id_xor_block(133) xor id_xor_block(135) xor id_xor_block(137) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(143) xor id_xor_block(145) xor id_xor_block(146) xor id_xor_block(148) xor id_xor_block(149) xor id_xor_block(150) xor id_xor_block(152) xor id_xor_block(155) xor id_xor_block(158) xor id_xor_block(159) xor id_xor_block(161) xor id_xor_block(163) xor id_xor_block(165) xor id_xor_block(166) xor id_xor_block(167) xor id_xor_block(168) xor id_xor_block(170) xor id_xor_block(171) xor id_xor_block(173) xor id_xor_block(176) xor id_xor_block(177) xor id_xor_block(179) xor id_xor_block(180) xor id_xor_block(182) xor id_xor_block(185) xor id_xor_block(189) xor id_xor_block(190) xor id_xor_block(191) xor id_xor_block(196) xor id_xor_block(197) xor id_xor_block(199) xor id_xor_block(200) xor id_xor_block(201) xor id_xor_block(202) xor id_xor_block(205) xor id_xor_block(207) xor id_xor_block(209) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(217) xor id_xor_block(221) xor id_xor_block(224) xor id_xor_block(225) xor id_xor_block(226) xor id_xor_block(227) xor id_xor_block(232) xor id_xor_block(234) xor id_xor_block(238) xor id_xor_block(239) xor id_xor_block(245);
	od_logic_block(6) <= id_xor_block(120) xor id_xor_block(121) xor id_xor_block(122) xor id_xor_block(123) xor id_xor_block(124) xor id_xor_block(127) xor id_xor_block(128) xor id_xor_block(131) xor id_xor_block(132) xor id_xor_block(133) xor id_xor_block(135) xor id_xor_block(138) xor id_xor_block(139) xor id_xor_block(140) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(143) xor id_xor_block(146) xor id_xor_block(147) xor id_xor_block(148) xor id_xor_block(151) xor id_xor_block(153) xor id_xor_block(154) xor id_xor_block(155) xor id_xor_block(162) xor id_xor_block(163) xor id_xor_block(165) xor id_xor_block(166) xor id_xor_block(169) xor id_xor_block(171) xor id_xor_block(173) xor id_xor_block(183) xor id_xor_block(185) xor id_xor_block(186) xor id_xor_block(187) xor id_xor_block(188) xor id_xor_block(189) xor id_xor_block(192) xor id_xor_block(193) xor id_xor_block(194) xor id_xor_block(195) xor id_xor_block(196) xor id_xor_block(199) xor id_xor_block(200) xor id_xor_block(203) xor id_xor_block(205) xor id_xor_block(208) xor id_xor_block(210) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(214) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(217) xor id_xor_block(219) xor id_xor_block(221) xor id_xor_block(222) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(228) xor id_xor_block(229) xor id_xor_block(230) xor id_xor_block(231) xor id_xor_block(232) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(235) xor id_xor_block(236) xor id_xor_block(237) xor id_xor_block(238) xor id_xor_block(246);
	od_logic_block(7) <= id_xor_block(121) xor id_xor_block(122) xor id_xor_block(123) xor id_xor_block(124) xor id_xor_block(125) xor id_xor_block(128) xor id_xor_block(129) xor id_xor_block(132) xor id_xor_block(133) xor id_xor_block(134) xor id_xor_block(136) xor id_xor_block(139) xor id_xor_block(140) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(143) xor id_xor_block(144) xor id_xor_block(147) xor id_xor_block(148) xor id_xor_block(149) xor id_xor_block(152) xor id_xor_block(154) xor id_xor_block(155) xor id_xor_block(156) xor id_xor_block(163) xor id_xor_block(164) xor id_xor_block(166) xor id_xor_block(167) xor id_xor_block(170) xor id_xor_block(172) xor id_xor_block(174) xor id_xor_block(184) xor id_xor_block(186) xor id_xor_block(187) xor id_xor_block(188) xor id_xor_block(189) xor id_xor_block(190) xor id_xor_block(193) xor id_xor_block(194) xor id_xor_block(195) xor id_xor_block(196) xor id_xor_block(197) xor id_xor_block(200) xor id_xor_block(201) xor id_xor_block(204) xor id_xor_block(206) xor id_xor_block(209) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(214) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(217) xor id_xor_block(218) xor id_xor_block(220) xor id_xor_block(222) xor id_xor_block(223) xor id_xor_block(224) xor id_xor_block(225) xor id_xor_block(229) xor id_xor_block(230) xor id_xor_block(231) xor id_xor_block(232) xor id_xor_block(233) xor id_xor_block(234) xor id_xor_block(235) xor id_xor_block(236) xor id_xor_block(237) xor id_xor_block(238) xor id_xor_block(239) xor id_xor_block(247);
	od_logic_block(8) <= id_xor_block(120) xor id_xor_block(121) xor id_xor_block(136) xor id_xor_block(137) xor id_xor_block(139) xor id_xor_block(153) xor id_xor_block(154) xor id_xor_block(157) xor id_xor_block(171) xor id_xor_block(172) xor id_xor_block(174) xor id_xor_block(175) xor id_xor_block(193) xor id_xor_block(206) xor id_xor_block(207) xor id_xor_block(210) xor id_xor_block(211) xor id_xor_block(227) xor id_xor_block(229) xor id_xor_block(248);
	od_logic_block(9) <= id_xor_block(121) xor id_xor_block(122) xor id_xor_block(137) xor id_xor_block(138) xor id_xor_block(140) xor id_xor_block(154) xor id_xor_block(155) xor id_xor_block(158) xor id_xor_block(172) xor id_xor_block(173) xor id_xor_block(175) xor id_xor_block(176) xor id_xor_block(194) xor id_xor_block(207) xor id_xor_block(208) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(228) xor id_xor_block(230) xor id_xor_block(249);
	od_logic_block(10) <= id_xor_block(122) xor id_xor_block(123) xor id_xor_block(138) xor id_xor_block(139) xor id_xor_block(141) xor id_xor_block(155) xor id_xor_block(156) xor id_xor_block(159) xor id_xor_block(173) xor id_xor_block(174) xor id_xor_block(176) xor id_xor_block(177) xor id_xor_block(195) xor id_xor_block(208) xor id_xor_block(209) xor id_xor_block(212) xor id_xor_block(213) xor id_xor_block(229) xor id_xor_block(231) xor id_xor_block(250);
	od_logic_block(11) <= id_xor_block(123) xor id_xor_block(124) xor id_xor_block(139) xor id_xor_block(140) xor id_xor_block(142) xor id_xor_block(156) xor id_xor_block(157) xor id_xor_block(160) xor id_xor_block(174) xor id_xor_block(175) xor id_xor_block(177) xor id_xor_block(178) xor id_xor_block(196) xor id_xor_block(209) xor id_xor_block(210) xor id_xor_block(213) xor id_xor_block(214) xor id_xor_block(230) xor id_xor_block(232) xor id_xor_block(251);
	od_logic_block(12) <= id_xor_block(124) xor id_xor_block(125) xor id_xor_block(140) xor id_xor_block(141) xor id_xor_block(143) xor id_xor_block(157) xor id_xor_block(158) xor id_xor_block(161) xor id_xor_block(175) xor id_xor_block(176) xor id_xor_block(178) xor id_xor_block(179) xor id_xor_block(197) xor id_xor_block(210) xor id_xor_block(211) xor id_xor_block(214) xor id_xor_block(215) xor id_xor_block(231) xor id_xor_block(233) xor id_xor_block(252);
	od_logic_block(13) <= id_xor_block(125) xor id_xor_block(126) xor id_xor_block(141) xor id_xor_block(142) xor id_xor_block(144) xor id_xor_block(158) xor id_xor_block(159) xor id_xor_block(162) xor id_xor_block(176) xor id_xor_block(177) xor id_xor_block(179) xor id_xor_block(180) xor id_xor_block(198) xor id_xor_block(211) xor id_xor_block(212) xor id_xor_block(215) xor id_xor_block(216) xor id_xor_block(232) xor id_xor_block(234) xor id_xor_block(253);
end rtl; 
